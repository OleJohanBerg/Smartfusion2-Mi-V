-- Version: 
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity MSS_025 is
	generic (
		INIT:std_logic_vector := x"0";
		ACT_UBITS:std_logic_vector := x"0";
		MEMORYFILE:string := "";
		RTC_MAIN_XTL_FREQ:real := 0.0;
		RTC_MAIN_XTL_MODE:string := "";
		DDR_CLK_FREQ:real := 0.0	);
   port( 
       CAN_RXBUS_MGPIO3A_H2F_A : out std_logic;
       CAN_RXBUS_MGPIO3A_H2F_B : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_A : out std_logic;
       CAN_TX_EBL_MGPIO4A_H2F_B : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_A : out std_logic;
       CAN_TXBUS_MGPIO2A_H2F_B : out std_logic;
       CLK_CONFIG_APB : out std_logic;
       COMMS_INT : out std_logic;
       CONFIG_PRESET_N : out std_logic;
       EDAC_ERROR : out std_logic_vector(7 downto 0);
       F_FM0_RDATA : out std_logic_vector(31 downto 0);
       F_FM0_READYOUT : out std_logic;
       F_FM0_RESP : out std_logic;
       F_HM0_ADDR : out std_logic_vector(31 downto 0);
       F_HM0_ENABLE : out std_logic;
       F_HM0_SEL : out std_logic;
       F_HM0_SIZE : out std_logic_vector(1 downto 0);
       F_HM0_TRANS1 : out std_logic;
       F_HM0_WDATA : out std_logic_vector(31 downto 0);
       F_HM0_WRITE : out std_logic;
       FAB_CHRGVBUS : out std_logic;
       FAB_DISCHRGVBUS : out std_logic;
       FAB_DMPULLDOWN : out std_logic;
       FAB_DPPULLDOWN : out std_logic;
       FAB_DRVVBUS : out std_logic;
       FAB_IDPULLUP : out std_logic;
       FAB_OPMODE : out std_logic_vector(1 downto 0);
       FAB_SUSPENDM : out std_logic;
       FAB_TERMSEL : out std_logic;
       FAB_TXVALID : out std_logic;
       FAB_VCONTROL : out std_logic_vector(3 downto 0);
       FAB_VCONTROLLOADM : out std_logic;
       FAB_XCVRSEL : out std_logic_vector(1 downto 0);
       FAB_XDATAOUT : out std_logic_vector(7 downto 0);
       FACC_GLMUX_SEL : out std_logic;
       FIC32_0_MASTER : out std_logic_vector(1 downto 0);
       FIC32_1_MASTER : out std_logic_vector(1 downto 0);
       FPGA_RESET_N : out std_logic;
       GTX_CLK : out std_logic;
       H2F_INTERRUPT : out std_logic_vector(15 downto 0);
       H2F_NMI : out std_logic;
       H2FCALIB : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_A : out std_logic;
       I2C0_SCL_MGPIO31B_H2F_B : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_A : out std_logic;
       I2C0_SDA_MGPIO30B_H2F_B : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_A : out std_logic;
       I2C1_SCL_MGPIO1A_H2F_B : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_A : out std_logic;
       I2C1_SDA_MGPIO0A_H2F_B : out std_logic;
       MDCF : out std_logic;
       MDOENF : out std_logic;
       MDOF : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_A : out std_logic;
       MMUART0_CTS_MGPIO19B_H2F_B : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_A : out std_logic;
       MMUART0_DCD_MGPIO22B_H2F_B : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_A : out std_logic;
       MMUART0_DSR_MGPIO20B_H2F_B : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_A : out std_logic;
       MMUART0_DTR_MGPIO18B_H2F_B : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_A : out std_logic;
       MMUART0_RI_MGPIO21B_H2F_B : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_A : out std_logic;
       MMUART0_RTS_MGPIO17B_H2F_B : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_A : out std_logic;
       MMUART0_RXD_MGPIO28B_H2F_B : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_A : out std_logic;
       MMUART0_SCK_MGPIO29B_H2F_B : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_A : out std_logic;
       MMUART0_TXD_MGPIO27B_H2F_B : out std_logic;
       MMUART1_DTR_MGPIO12B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_A : out std_logic;
       MMUART1_RTS_MGPIO11B_H2F_B : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_A : out std_logic;
       MMUART1_RXD_MGPIO26B_H2F_B : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_A : out std_logic;
       MMUART1_SCK_MGPIO25B_H2F_B : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_A : out std_logic;
       MMUART1_TXD_MGPIO24B_H2F_B : out std_logic;
       MPLL_LOCK : out std_logic;
       PER2_FABRIC_PADDR : out std_logic_vector(15 downto 2);
       PER2_FABRIC_PENABLE : out std_logic;
       PER2_FABRIC_PSEL : out std_logic;
       PER2_FABRIC_PWDATA : out std_logic_vector(31 downto 0);
       PER2_FABRIC_PWRITE : out std_logic;
       RTC_MATCH : out std_logic;
       SLEEPDEEP : out std_logic;
       SLEEPHOLDACK : out std_logic;
       SLEEPING : out std_logic;
       SMBALERT_NO0 : out std_logic;
       SMBALERT_NO1 : out std_logic;
       SMBSUS_NO0 : out std_logic;
       SMBSUS_NO1 : out std_logic;
       SPI0_CLK_OUT : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_A : out std_logic;
       SPI0_SDI_MGPIO5A_H2F_B : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_A : out std_logic;
       SPI0_SDO_MGPIO6A_H2F_B : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_A : out std_logic;
       SPI0_SS0_MGPIO7A_H2F_B : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_A : out std_logic;
       SPI0_SS1_MGPIO8A_H2F_B : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_A : out std_logic;
       SPI0_SS2_MGPIO9A_H2F_B : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_A : out std_logic;
       SPI0_SS3_MGPIO10A_H2F_B : out std_logic;
       SPI0_SS4_MGPIO19A_H2F_A : out std_logic;
       SPI0_SS5_MGPIO20A_H2F_A : out std_logic;
       SPI0_SS6_MGPIO21A_H2F_A : out std_logic;
       SPI0_SS7_MGPIO22A_H2F_A : out std_logic;
       SPI1_CLK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_A : out std_logic;
       SPI1_SDI_MGPIO11A_H2F_B : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_A : out std_logic;
       SPI1_SDO_MGPIO12A_H2F_B : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_A : out std_logic;
       SPI1_SS0_MGPIO13A_H2F_B : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_A : out std_logic;
       SPI1_SS1_MGPIO14A_H2F_B : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_A : out std_logic;
       SPI1_SS2_MGPIO15A_H2F_B : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_A : out std_logic;
       SPI1_SS3_MGPIO16A_H2F_B : out std_logic;
       SPI1_SS4_MGPIO17A_H2F_A : out std_logic;
       SPI1_SS5_MGPIO18A_H2F_A : out std_logic;
       SPI1_SS6_MGPIO23A_H2F_A : out std_logic;
       SPI1_SS7_MGPIO24A_H2F_A : out std_logic;
       TCGF : out std_logic_vector(9 downto 0);
       TRACECLK : out std_logic;
       TRACEDATA : out std_logic_vector(3 downto 0);
       TX_CLK : out std_logic;
       TX_ENF : out std_logic;
       TX_ERRF : out std_logic;
       TXCTL_EN_RIF : out std_logic;
       TXD_RIF : out std_logic_vector(3 downto 0);
       TXDF : out std_logic_vector(7 downto 0);
       TXEV : out std_logic;
       WDOGTIMEOUT : out std_logic;
       F_ARREADY_HREADYOUT1 : out std_logic;
       F_AWREADY_HREADYOUT0 : out std_logic;
       F_BID : out std_logic_vector(3 downto 0);
       F_BRESP_HRESP0 : out std_logic_vector(1 downto 0);
       F_BVALID : out std_logic;
       F_RDATA_HRDATA01 : out std_logic_vector(63 downto 0);
       F_RID : out std_logic_vector(3 downto 0);
       F_RLAST : out std_logic;
       F_RRESP_HRESP1 : out std_logic_vector(1 downto 0);
       F_RVALID : out std_logic;
       F_WREADY : out std_logic;
       MDDR_FABRIC_PRDATA : out std_logic_vector(15 downto 0);
       MDDR_FABRIC_PREADY : out std_logic;
       MDDR_FABRIC_PSLVERR : out std_logic;
       CAN_RXBUS_F2H_SCP : in std_logic;
       CAN_TX_EBL_F2H_SCP : in std_logic;
       CAN_TXBUS_F2H_SCP : in std_logic;
       COLF : in std_logic;
       CRSF : in std_logic;
       F2_DMAREADY : in std_logic_vector(1 downto 0);
       F2H_INTERRUPT : in std_logic_vector(15 downto 0);
       F2HCALIB : in std_logic;
       F_DMAREADY : in std_logic_vector(1 downto 0);
       F_FM0_ADDR : in std_logic_vector(31 downto 0);
       F_FM0_ENABLE : in std_logic;
       F_FM0_MASTLOCK : in std_logic;
       F_FM0_READY : in std_logic;
       F_FM0_SEL : in std_logic;
       F_FM0_SIZE : in std_logic_vector(1 downto 0);
       F_FM0_TRANS1 : in std_logic;
       F_FM0_WDATA : in std_logic_vector(31 downto 0);
       F_FM0_WRITE : in std_logic;
       F_HM0_RDATA : in std_logic_vector(31 downto 0);
       F_HM0_READY : in std_logic;
       F_HM0_RESP : in std_logic;
       FAB_AVALID : in std_logic;
       FAB_HOSTDISCON : in std_logic;
       FAB_IDDIG : in std_logic;
       FAB_LINESTATE : in std_logic_vector(1 downto 0);
       FAB_M3_RESET_N : in std_logic;
       FAB_PLL_LOCK : in std_logic;
       FAB_RXACTIVE : in std_logic;
       FAB_RXERROR : in std_logic;
       FAB_RXVALID : in std_logic;
       FAB_RXVALIDH : in std_logic;
       FAB_SESSEND : in std_logic;
       FAB_TXREADY : in std_logic;
       FAB_VBUSVALID : in std_logic;
       FAB_VSTATUS : in std_logic_vector(7 downto 0);
       FAB_XDATAIN : in std_logic_vector(7 downto 0);
       GTX_CLKPF : in std_logic;
       I2C0_BCLK : in std_logic;
       I2C0_SCL_F2H_SCP : in std_logic;
       I2C0_SDA_F2H_SCP : in std_logic;
       I2C1_BCLK : in std_logic;
       I2C1_SCL_F2H_SCP : in std_logic;
       I2C1_SDA_F2H_SCP : in std_logic;
       MDIF : in std_logic;
       MGPIO0A_F2H_GPIN : in std_logic;
       MGPIO10A_F2H_GPIN : in std_logic;
       MGPIO11A_F2H_GPIN : in std_logic;
       MGPIO11B_F2H_GPIN : in std_logic;
       MGPIO12A_F2H_GPIN : in std_logic;
       MGPIO13A_F2H_GPIN : in std_logic;
       MGPIO14A_F2H_GPIN : in std_logic;
       MGPIO15A_F2H_GPIN : in std_logic;
       MGPIO16A_F2H_GPIN : in std_logic;
       MGPIO17B_F2H_GPIN : in std_logic;
       MGPIO18B_F2H_GPIN : in std_logic;
       MGPIO19B_F2H_GPIN : in std_logic;
       MGPIO1A_F2H_GPIN : in std_logic;
       MGPIO20B_F2H_GPIN : in std_logic;
       MGPIO21B_F2H_GPIN : in std_logic;
       MGPIO22B_F2H_GPIN : in std_logic;
       MGPIO24B_F2H_GPIN : in std_logic;
       MGPIO25B_F2H_GPIN : in std_logic;
       MGPIO26B_F2H_GPIN : in std_logic;
       MGPIO27B_F2H_GPIN : in std_logic;
       MGPIO28B_F2H_GPIN : in std_logic;
       MGPIO29B_F2H_GPIN : in std_logic;
       MGPIO2A_F2H_GPIN : in std_logic;
       MGPIO30B_F2H_GPIN : in std_logic;
       MGPIO31B_F2H_GPIN : in std_logic;
       MGPIO3A_F2H_GPIN : in std_logic;
       MGPIO4A_F2H_GPIN : in std_logic;
       MGPIO5A_F2H_GPIN : in std_logic;
       MGPIO6A_F2H_GPIN : in std_logic;
       MGPIO7A_F2H_GPIN : in std_logic;
       MGPIO8A_F2H_GPIN : in std_logic;
       MGPIO9A_F2H_GPIN : in std_logic;
       MMUART0_CTS_F2H_SCP : in std_logic;
       MMUART0_DCD_F2H_SCP : in std_logic;
       MMUART0_DSR_F2H_SCP : in std_logic;
       MMUART0_DTR_F2H_SCP : in std_logic;
       MMUART0_RI_F2H_SCP : in std_logic;
       MMUART0_RTS_F2H_SCP : in std_logic;
       MMUART0_RXD_F2H_SCP : in std_logic;
       MMUART0_SCK_F2H_SCP : in std_logic;
       MMUART0_TXD_F2H_SCP : in std_logic;
       MMUART1_CTS_F2H_SCP : in std_logic;
       MMUART1_DCD_F2H_SCP : in std_logic;
       MMUART1_DSR_F2H_SCP : in std_logic;
       MMUART1_RI_F2H_SCP : in std_logic;
       MMUART1_RTS_F2H_SCP : in std_logic;
       MMUART1_RXD_F2H_SCP : in std_logic;
       MMUART1_SCK_F2H_SCP : in std_logic;
       MMUART1_TXD_F2H_SCP : in std_logic;
       PER2_FABRIC_PRDATA : in std_logic_vector(31 downto 0);
       PER2_FABRIC_PREADY : in std_logic;
       PER2_FABRIC_PSLVERR : in std_logic;
       RCGF : in std_logic_vector(9 downto 0);
       RX_CLKPF : in std_logic;
       RX_DVF : in std_logic;
       RX_ERRF : in std_logic;
       RX_EV : in std_logic;
       RXDF : in std_logic_vector(7 downto 0);
       SLEEPHOLDREQ : in std_logic;
       SMBALERT_NI0 : in std_logic;
       SMBALERT_NI1 : in std_logic;
       SMBSUS_NI0 : in std_logic;
       SMBSUS_NI1 : in std_logic;
       SPI0_CLK_IN : in std_logic;
       SPI0_SDI_F2H_SCP : in std_logic;
       SPI0_SDO_F2H_SCP : in std_logic;
       SPI0_SS0_F2H_SCP : in std_logic;
       SPI0_SS1_F2H_SCP : in std_logic;
       SPI0_SS2_F2H_SCP : in std_logic;
       SPI0_SS3_F2H_SCP : in std_logic;
       SPI1_CLK_IN : in std_logic;
       SPI1_SDI_F2H_SCP : in std_logic;
       SPI1_SDO_F2H_SCP : in std_logic;
       SPI1_SS0_F2H_SCP : in std_logic;
       SPI1_SS1_F2H_SCP : in std_logic;
       SPI1_SS2_F2H_SCP : in std_logic;
       SPI1_SS3_F2H_SCP : in std_logic;
       TX_CLKPF : in std_logic;
       USER_MSS_GPIO_RESET_N : in std_logic;
       USER_MSS_RESET_N : in std_logic;
       XCLK_FAB : in std_logic;
       CLK_BASE : in std_logic;
       CLK_MDDR_APB : in std_logic;
       F_ARADDR_HADDR1 : in std_logic_vector(31 downto 0);
       F_ARBURST_HTRANS1 : in std_logic_vector(1 downto 0);
       F_ARID_HSEL1 : in std_logic_vector(3 downto 0);
       F_ARLEN_HBURST1 : in std_logic_vector(3 downto 0);
       F_ARLOCK_HMASTLOCK1 : in std_logic_vector(1 downto 0);
       F_ARSIZE_HSIZE1 : in std_logic_vector(1 downto 0);
       F_ARVALID_HWRITE1 : in std_logic;
       F_AWADDR_HADDR0 : in std_logic_vector(31 downto 0);
       F_AWBURST_HTRANS0 : in std_logic_vector(1 downto 0);
       F_AWID_HSEL0 : in std_logic_vector(3 downto 0);
       F_AWLEN_HBURST0 : in std_logic_vector(3 downto 0);
       F_AWLOCK_HMASTLOCK0 : in std_logic_vector(1 downto 0);
       F_AWSIZE_HSIZE0 : in std_logic_vector(1 downto 0);
       F_AWVALID_HWRITE0 : in std_logic;
       F_BREADY : in std_logic;
       F_RMW_AXI : in std_logic;
       F_RREADY : in std_logic;
       F_WDATA_HWDATA01 : in std_logic_vector(63 downto 0);
       F_WID_HREADY01 : in std_logic_vector(3 downto 0);
       F_WLAST : in std_logic;
       F_WSTRB : in std_logic_vector(7 downto 0);
       F_WVALID : in std_logic;
       FPGA_MDDR_ARESET_N : in std_logic;
       MDDR_FABRIC_PADDR : in std_logic_vector(10 downto 2);
       MDDR_FABRIC_PENABLE : in std_logic;
       MDDR_FABRIC_PSEL : in std_logic;
       MDDR_FABRIC_PWDATA : in std_logic_vector(15 downto 0);
       MDDR_FABRIC_PWRITE : in std_logic;
       PRESET_N : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN : in std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN : in std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN : in std_logic;
       DM_IN : in std_logic_vector(2 downto 0);
       DRAM_DQ_IN : in std_logic_vector(17 downto 0);
       DRAM_DQS_IN : in std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_IN : in std_logic_vector(1 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN : in std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN : in std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN : in std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN : in std_logic;
       MGPIO25A_IN : in std_logic;
       MGPIO26A_IN : in std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN : in std_logic;
       MMUART0_DCD_MGPIO22B_IN : in std_logic;
       MMUART0_DSR_MGPIO20B_IN : in std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN : in std_logic;
       MMUART0_RI_MGPIO21B_IN : in std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN : in std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_IN : in std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN : in std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN : in std_logic;
       MMUART1_CTS_MGPIO13B_IN : in std_logic;
       MMUART1_DCD_MGPIO16B_IN : in std_logic;
       MMUART1_DSR_MGPIO14B_IN : in std_logic;
       MMUART1_DTR_MGPIO12B_IN : in std_logic;
       MMUART1_RI_MGPIO15B_IN : in std_logic;
       MMUART1_RTS_MGPIO11B_IN : in std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN : in std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN : in std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN : in std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN : in std_logic;
       RGMII_MDC_RMII_MDC_IN : in std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN : in std_logic;
       RGMII_RX_CLK_IN : in std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN : in std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN : in std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN : in std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN : in std_logic;
       RGMII_RXD3_USBB_DATA4_IN : in std_logic;
       RGMII_TX_CLK_IN : in std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN : in std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN : in std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN : in std_logic;
       RGMII_TXD2_USBB_DATA5_IN : in std_logic;
       RGMII_TXD3_USBB_DATA6_IN : in std_logic;
       SPI0_SCK_USBA_XCLK_IN : in std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_IN : in std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_IN : in std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_IN : in std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN : in std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN : in std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN : in std_logic;
       SPI0_SS4_MGPIO19A_IN : in std_logic;
       SPI0_SS5_MGPIO20A_IN : in std_logic;
       SPI0_SS6_MGPIO21A_IN : in std_logic;
       SPI0_SS7_MGPIO22A_IN : in std_logic;
       SPI1_SCK_IN : in std_logic;
       SPI1_SDI_MGPIO11A_IN : in std_logic;
       SPI1_SDO_MGPIO12A_IN : in std_logic;
       SPI1_SS0_MGPIO13A_IN : in std_logic;
       SPI1_SS1_MGPIO14A_IN : in std_logic;
       SPI1_SS2_MGPIO15A_IN : in std_logic;
       SPI1_SS3_MGPIO16A_IN : in std_logic;
       SPI1_SS4_MGPIO17A_IN : in std_logic;
       SPI1_SS5_MGPIO18A_IN : in std_logic;
       SPI1_SS6_MGPIO23A_IN : in std_logic;
       SPI1_SS7_MGPIO24A_IN : in std_logic;
       USBC_XCLK_IN : in std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT : out std_logic;
       DRAM_ADDR : out std_logic_vector(15 downto 0);
       DRAM_BA : out std_logic_vector(2 downto 0);
       DRAM_CASN : out std_logic;
       DRAM_CKE : out std_logic;
       DRAM_CLK : out std_logic;
       DRAM_CSN : out std_logic;
       DRAM_DM_RDQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_DQ_OUT : out std_logic_vector(17 downto 0);
       DRAM_DQS_OUT : out std_logic_vector(2 downto 0);
       DRAM_FIFO_WE_OUT : out std_logic_vector(1 downto 0);
       DRAM_ODT : out std_logic;
       DRAM_RASN : out std_logic;
       DRAM_RSTN : out std_logic;
       DRAM_WEN : out std_logic;
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT : out std_logic;
       MGPIO25A_OUT : out std_logic;
       MGPIO26A_OUT : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT : out std_logic;
       MMUART0_DCD_MGPIO22B_OUT : out std_logic;
       MMUART0_DSR_MGPIO20B_OUT : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT : out std_logic;
       MMUART0_RI_MGPIO21B_OUT : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT : out std_logic;
       MMUART1_CTS_MGPIO13B_OUT : out std_logic;
       MMUART1_DCD_MGPIO16B_OUT : out std_logic;
       MMUART1_DSR_MGPIO14B_OUT : out std_logic;
       MMUART1_DTR_MGPIO12B_OUT : out std_logic;
       MMUART1_RI_MGPIO15B_OUT : out std_logic;
       MMUART1_RTS_MGPIO11B_OUT : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT : out std_logic;
       RGMII_MDC_RMII_MDC_OUT : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT : out std_logic;
       RGMII_RX_CLK_OUT : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT : out std_logic;
       RGMII_RXD3_USBB_DATA4_OUT : out std_logic;
       RGMII_TX_CLK_OUT : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT : out std_logic;
       RGMII_TXD2_USBB_DATA5_OUT : out std_logic;
       RGMII_TXD3_USBB_DATA6_OUT : out std_logic;
       SPI0_SCK_USBA_XCLK_OUT : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OUT : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT : out std_logic;
       SPI0_SS4_MGPIO19A_OUT : out std_logic;
       SPI0_SS5_MGPIO20A_OUT : out std_logic;
       SPI0_SS6_MGPIO21A_OUT : out std_logic;
       SPI0_SS7_MGPIO22A_OUT : out std_logic;
       SPI1_SCK_OUT : out std_logic;
       SPI1_SDI_MGPIO11A_OUT : out std_logic;
       SPI1_SDO_MGPIO12A_OUT : out std_logic;
       SPI1_SS0_MGPIO13A_OUT : out std_logic;
       SPI1_SS1_MGPIO14A_OUT : out std_logic;
       SPI1_SS2_MGPIO15A_OUT : out std_logic;
       SPI1_SS3_MGPIO16A_OUT : out std_logic;
       SPI1_SS4_MGPIO17A_OUT : out std_logic;
       SPI1_SS5_MGPIO18A_OUT : out std_logic;
       SPI1_SS6_MGPIO23A_OUT : out std_logic;
       SPI1_SS7_MGPIO24A_OUT : out std_logic;
       USBC_XCLK_OUT : out std_logic;
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE : out std_logic;
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE : out std_logic;
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE : out std_logic;
       DM_OE : out std_logic_vector(2 downto 0);
       DRAM_DQ_OE : out std_logic_vector(17 downto 0);
       DRAM_DQS_OE : out std_logic_vector(2 downto 0);
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE : out std_logic;
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE : out std_logic;
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE : out std_logic;
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE : out std_logic;
       MGPIO25A_OE : out std_logic;
       MGPIO26A_OE : out std_logic;
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE : out std_logic;
       MMUART0_DCD_MGPIO22B_OE : out std_logic;
       MMUART0_DSR_MGPIO20B_OE : out std_logic;
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE : out std_logic;
       MMUART0_RI_MGPIO21B_OE : out std_logic;
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE : out std_logic;
       MMUART0_RXD_USBC_STP_MGPIO28B_OE : out std_logic;
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE : out std_logic;
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE : out std_logic;
       MMUART1_CTS_MGPIO13B_OE : out std_logic;
       MMUART1_DCD_MGPIO16B_OE : out std_logic;
       MMUART1_DSR_MGPIO14B_OE : out std_logic;
       MMUART1_DTR_MGPIO12B_OE : out std_logic;
       MMUART1_RI_MGPIO15B_OE : out std_logic;
       MMUART1_RTS_MGPIO11B_OE : out std_logic;
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE : out std_logic;
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE : out std_logic;
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE : out std_logic;
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE : out std_logic;
       RGMII_MDC_RMII_MDC_OE : out std_logic;
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE : out std_logic;
       RGMII_RX_CLK_OE : out std_logic;
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE : out std_logic;
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE : out std_logic;
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE : out std_logic;
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE : out std_logic;
       RGMII_RXD3_USBB_DATA4_OE : out std_logic;
       RGMII_TX_CLK_OE : out std_logic;
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE : out std_logic;
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE : out std_logic;
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE : out std_logic;
       RGMII_TXD2_USBB_DATA5_OE : out std_logic;
       RGMII_TXD3_USBB_DATA6_OE : out std_logic;
       SPI0_SCK_USBA_XCLK_OE : out std_logic;
       SPI0_SDI_USBA_DIR_MGPIO5A_OE : out std_logic;
       SPI0_SDO_USBA_STP_MGPIO6A_OE : out std_logic;
       SPI0_SS0_USBA_NXT_MGPIO7A_OE : out std_logic;
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE : out std_logic;
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE : out std_logic;
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE : out std_logic;
       SPI0_SS4_MGPIO19A_OE : out std_logic;
       SPI0_SS5_MGPIO20A_OE : out std_logic;
       SPI0_SS6_MGPIO21A_OE : out std_logic;
       SPI0_SS7_MGPIO22A_OE : out std_logic;
       SPI1_SCK_OE : out std_logic;
       SPI1_SDI_MGPIO11A_OE : out std_logic;
       SPI1_SDO_MGPIO12A_OE : out std_logic;
       SPI1_SS0_MGPIO13A_OE : out std_logic;
       SPI1_SS1_MGPIO14A_OE : out std_logic;
       SPI1_SS2_MGPIO15A_OE : out std_logic;
       SPI1_SS3_MGPIO16A_OE : out std_logic;
       SPI1_SS4_MGPIO17A_OE : out std_logic;
       SPI1_SS5_MGPIO18A_OE : out std_logic;
       SPI1_SS6_MGPIO23A_OE : out std_logic;
       SPI1_SS7_MGPIO24A_OE : out std_logic;
       USBC_XCLK_OE : out std_logic
   );
end MSS_025;
architecture DEF_ARCH of MSS_025 is 

   attribute black_box : boolean;
   attribute black_box of DEF_ARCH : architecture is true;
   attribute ment_tsu0: string;
   attribute ment_tsu0 of DEF_ARCH : architecture is " CAN_RXBUS_F2H_SCP->CLK_BASE=1.470";
   attribute ment_tsu1: string;
   attribute ment_tsu1 of DEF_ARCH : architecture is " F2HCALIB->CLK_BASE=1.317";
   attribute ment_tsu2: string;
   attribute ment_tsu2 of DEF_ARCH : architecture is " F2H_INTERRUPT[0]->CLK_BASE=0.961";
   attribute ment_tsu3: string;
   attribute ment_tsu3 of DEF_ARCH : architecture is " F2H_INTERRUPT[10]->CLK_BASE=1.091";
   attribute ment_tsu4: string;
   attribute ment_tsu4 of DEF_ARCH : architecture is " F2H_INTERRUPT[11]->CLK_BASE=1.027";
   attribute ment_tsu5: string;
   attribute ment_tsu5 of DEF_ARCH : architecture is " F2H_INTERRUPT[12]->CLK_BASE=1.013";
   attribute ment_tsu6: string;
   attribute ment_tsu6 of DEF_ARCH : architecture is " F2H_INTERRUPT[13]->CLK_BASE=0.996";
   attribute ment_tsu7: string;
   attribute ment_tsu7 of DEF_ARCH : architecture is " F2H_INTERRUPT[14]->CLK_BASE=1.027";
   attribute ment_tsu8: string;
   attribute ment_tsu8 of DEF_ARCH : architecture is " F2H_INTERRUPT[15]->CLK_BASE=0.999";
   attribute ment_tsu9: string;
   attribute ment_tsu9 of DEF_ARCH : architecture is " F2H_INTERRUPT[1]->CLK_BASE=0.968";
   attribute ment_tsu10: string;
   attribute ment_tsu10 of DEF_ARCH : architecture is " F2H_INTERRUPT[2]->CLK_BASE=1.029";
   attribute ment_tsu11: string;
   attribute ment_tsu11 of DEF_ARCH : architecture is " F2H_INTERRUPT[3]->CLK_BASE=0.962";
   attribute ment_tsu12: string;
   attribute ment_tsu12 of DEF_ARCH : architecture is " F2H_INTERRUPT[4]->CLK_BASE=1.009";
   attribute ment_tsu13: string;
   attribute ment_tsu13 of DEF_ARCH : architecture is " F2H_INTERRUPT[5]->CLK_BASE=1.048";
   attribute ment_tsu14: string;
   attribute ment_tsu14 of DEF_ARCH : architecture is " F2H_INTERRUPT[6]->CLK_BASE=0.999";
   attribute ment_tsu15: string;
   attribute ment_tsu15 of DEF_ARCH : architecture is " F2H_INTERRUPT[7]->CLK_BASE=0.994";
   attribute ment_tsu16: string;
   attribute ment_tsu16 of DEF_ARCH : architecture is " F2H_INTERRUPT[8]->CLK_BASE=1.030";
   attribute ment_tsu17: string;
   attribute ment_tsu17 of DEF_ARCH : architecture is " F2H_INTERRUPT[9]->CLK_BASE=0.985";
   attribute ment_tsu18: string;
   attribute ment_tsu18 of DEF_ARCH : architecture is " F_FM0_ADDR[0]->CLK_BASE=0.966";
   attribute ment_tsu19: string;
   attribute ment_tsu19 of DEF_ARCH : architecture is " F_FM0_ADDR[10]->CLK_BASE=0.996";
   attribute ment_tsu20: string;
   attribute ment_tsu20 of DEF_ARCH : architecture is " F_FM0_ADDR[11]->CLK_BASE=1.020";
   attribute ment_tsu21: string;
   attribute ment_tsu21 of DEF_ARCH : architecture is " F_FM0_ADDR[12]->CLK_BASE=1.051";
   attribute ment_tsu22: string;
   attribute ment_tsu22 of DEF_ARCH : architecture is " F_FM0_ADDR[13]->CLK_BASE=1.148";
   attribute ment_tsu23: string;
   attribute ment_tsu23 of DEF_ARCH : architecture is " F_FM0_ADDR[14]->CLK_BASE=1.033";
   attribute ment_tsu24: string;
   attribute ment_tsu24 of DEF_ARCH : architecture is " F_FM0_ADDR[15]->CLK_BASE=1.147";
   attribute ment_tsu25: string;
   attribute ment_tsu25 of DEF_ARCH : architecture is " F_FM0_ADDR[16]->CLK_BASE=1.022";
   attribute ment_tsu26: string;
   attribute ment_tsu26 of DEF_ARCH : architecture is " F_FM0_ADDR[17]->CLK_BASE=0.593";
   attribute ment_tsu27: string;
   attribute ment_tsu27 of DEF_ARCH : architecture is " F_FM0_ADDR[18]->CLK_BASE=0.782";
   attribute ment_tsu28: string;
   attribute ment_tsu28 of DEF_ARCH : architecture is " F_FM0_ADDR[19]->CLK_BASE=0.567";
   attribute ment_tsu29: string;
   attribute ment_tsu29 of DEF_ARCH : architecture is " F_FM0_ADDR[1]->CLK_BASE=0.987";
   attribute ment_tsu30: string;
   attribute ment_tsu30 of DEF_ARCH : architecture is " F_FM0_ADDR[20]->CLK_BASE=0.589";
   attribute ment_tsu31: string;
   attribute ment_tsu31 of DEF_ARCH : architecture is " F_FM0_ADDR[21]->CLK_BASE=0.540";
   attribute ment_tsu32: string;
   attribute ment_tsu32 of DEF_ARCH : architecture is " F_FM0_ADDR[22]->CLK_BASE=0.586";
   attribute ment_tsu33: string;
   attribute ment_tsu33 of DEF_ARCH : architecture is " F_FM0_ADDR[23]->CLK_BASE=0.601";
   attribute ment_tsu34: string;
   attribute ment_tsu34 of DEF_ARCH : architecture is " F_FM0_ADDR[24]->CLK_BASE=0.595";
   attribute ment_tsu35: string;
   attribute ment_tsu35 of DEF_ARCH : architecture is " F_FM0_ADDR[25]->CLK_BASE=0.685";
   attribute ment_tsu36: string;
   attribute ment_tsu36 of DEF_ARCH : architecture is " F_FM0_ADDR[26]->CLK_BASE=0.727";
   attribute ment_tsu37: string;
   attribute ment_tsu37 of DEF_ARCH : architecture is " F_FM0_ADDR[27]->CLK_BASE=0.742";
   attribute ment_tsu38: string;
   attribute ment_tsu38 of DEF_ARCH : architecture is " F_FM0_ADDR[28]->CLK_BASE=0.736";
   attribute ment_tsu39: string;
   attribute ment_tsu39 of DEF_ARCH : architecture is " F_FM0_ADDR[29]->CLK_BASE=0.558";
   attribute ment_tsu40: string;
   attribute ment_tsu40 of DEF_ARCH : architecture is " F_FM0_ADDR[2]->CLK_BASE=0.398";
   attribute ment_tsu41: string;
   attribute ment_tsu41 of DEF_ARCH : architecture is " F_FM0_ADDR[30]->CLK_BASE=0.660";
   attribute ment_tsu42: string;
   attribute ment_tsu42 of DEF_ARCH : architecture is " F_FM0_ADDR[31]->CLK_BASE=0.579";
   attribute ment_tsu43: string;
   attribute ment_tsu43 of DEF_ARCH : architecture is " F_FM0_ADDR[3]->CLK_BASE=1.001";
   attribute ment_tsu44: string;
   attribute ment_tsu44 of DEF_ARCH : architecture is " F_FM0_ADDR[4]->CLK_BASE=1.004";
   attribute ment_tsu45: string;
   attribute ment_tsu45 of DEF_ARCH : architecture is " F_FM0_ADDR[5]->CLK_BASE=0.934";
   attribute ment_tsu46: string;
   attribute ment_tsu46 of DEF_ARCH : architecture is " F_FM0_ADDR[6]->CLK_BASE=0.984";
   attribute ment_tsu47: string;
   attribute ment_tsu47 of DEF_ARCH : architecture is " F_FM0_ADDR[7]->CLK_BASE=1.006";
   attribute ment_tsu48: string;
   attribute ment_tsu48 of DEF_ARCH : architecture is " F_FM0_ADDR[8]->CLK_BASE=1.021";
   attribute ment_tsu49: string;
   attribute ment_tsu49 of DEF_ARCH : architecture is " F_FM0_ADDR[9]->CLK_BASE=1.048";
   attribute ment_tsu50: string;
   attribute ment_tsu50 of DEF_ARCH : architecture is " F_FM0_MASTLOCK->CLK_BASE=0.564";
   attribute ment_tsu51: string;
   attribute ment_tsu51 of DEF_ARCH : architecture is " F_FM0_READY->CLK_BASE=0.698";
   attribute ment_tsu52: string;
   attribute ment_tsu52 of DEF_ARCH : architecture is " F_FM0_SEL->CLK_BASE=1.125";
   attribute ment_tsu53: string;
   attribute ment_tsu53 of DEF_ARCH : architecture is " F_FM0_SIZE[0]->CLK_BASE=0.381";
   attribute ment_tsu54: string;
   attribute ment_tsu54 of DEF_ARCH : architecture is " F_FM0_SIZE[1]->CLK_BASE=0.438";
   attribute ment_tsu55: string;
   attribute ment_tsu55 of DEF_ARCH : architecture is " F_FM0_TRANS1->CLK_BASE=0.726";
   attribute ment_tsu56: string;
   attribute ment_tsu56 of DEF_ARCH : architecture is " F_FM0_WDATA[0]->CLK_BASE=0.493";
   attribute ment_tsu57: string;
   attribute ment_tsu57 of DEF_ARCH : architecture is " F_FM0_WDATA[10]->CLK_BASE=0.361";
   attribute ment_tsu58: string;
   attribute ment_tsu58 of DEF_ARCH : architecture is " F_FM0_WDATA[11]->CLK_BASE=0.393";
   attribute ment_tsu59: string;
   attribute ment_tsu59 of DEF_ARCH : architecture is " F_FM0_WDATA[12]->CLK_BASE=0.404";
   attribute ment_tsu60: string;
   attribute ment_tsu60 of DEF_ARCH : architecture is " F_FM0_WDATA[13]->CLK_BASE=0.477";
   attribute ment_tsu61: string;
   attribute ment_tsu61 of DEF_ARCH : architecture is " F_FM0_WDATA[14]->CLK_BASE=0.670";
   attribute ment_tsu62: string;
   attribute ment_tsu62 of DEF_ARCH : architecture is " F_FM0_WDATA[15]->CLK_BASE=0.432";
   attribute ment_tsu63: string;
   attribute ment_tsu63 of DEF_ARCH : architecture is " F_FM0_WDATA[16]->CLK_BASE=0.425";
   attribute ment_tsu64: string;
   attribute ment_tsu64 of DEF_ARCH : architecture is " F_FM0_WDATA[17]->CLK_BASE=0.554";
   attribute ment_tsu65: string;
   attribute ment_tsu65 of DEF_ARCH : architecture is " F_FM0_WDATA[18]->CLK_BASE=0.546";
   attribute ment_tsu66: string;
   attribute ment_tsu66 of DEF_ARCH : architecture is " F_FM0_WDATA[19]->CLK_BASE=0.381";
   attribute ment_tsu67: string;
   attribute ment_tsu67 of DEF_ARCH : architecture is " F_FM0_WDATA[1]->CLK_BASE=0.452";
   attribute ment_tsu68: string;
   attribute ment_tsu68 of DEF_ARCH : architecture is " F_FM0_WDATA[20]->CLK_BASE=0.399";
   attribute ment_tsu69: string;
   attribute ment_tsu69 of DEF_ARCH : architecture is " F_FM0_WDATA[21]->CLK_BASE=0.388";
   attribute ment_tsu70: string;
   attribute ment_tsu70 of DEF_ARCH : architecture is " F_FM0_WDATA[22]->CLK_BASE=0.443";
   attribute ment_tsu71: string;
   attribute ment_tsu71 of DEF_ARCH : architecture is " F_FM0_WDATA[23]->CLK_BASE=0.355";
   attribute ment_tsu72: string;
   attribute ment_tsu72 of DEF_ARCH : architecture is " F_FM0_WDATA[24]->CLK_BASE=0.486";
   attribute ment_tsu73: string;
   attribute ment_tsu73 of DEF_ARCH : architecture is " F_FM0_WDATA[25]->CLK_BASE=0.402";
   attribute ment_tsu74: string;
   attribute ment_tsu74 of DEF_ARCH : architecture is " F_FM0_WDATA[26]->CLK_BASE=0.396";
   attribute ment_tsu75: string;
   attribute ment_tsu75 of DEF_ARCH : architecture is " F_FM0_WDATA[27]->CLK_BASE=0.465";
   attribute ment_tsu76: string;
   attribute ment_tsu76 of DEF_ARCH : architecture is " F_FM0_WDATA[28]->CLK_BASE=0.418";
   attribute ment_tsu77: string;
   attribute ment_tsu77 of DEF_ARCH : architecture is " F_FM0_WDATA[29]->CLK_BASE=0.383";
   attribute ment_tsu78: string;
   attribute ment_tsu78 of DEF_ARCH : architecture is " F_FM0_WDATA[2]->CLK_BASE=0.388";
   attribute ment_tsu79: string;
   attribute ment_tsu79 of DEF_ARCH : architecture is " F_FM0_WDATA[30]->CLK_BASE=0.359";
   attribute ment_tsu80: string;
   attribute ment_tsu80 of DEF_ARCH : architecture is " F_FM0_WDATA[31]->CLK_BASE=0.365";
   attribute ment_tsu81: string;
   attribute ment_tsu81 of DEF_ARCH : architecture is " F_FM0_WDATA[3]->CLK_BASE=0.387";
   attribute ment_tsu82: string;
   attribute ment_tsu82 of DEF_ARCH : architecture is " F_FM0_WDATA[4]->CLK_BASE=0.403";
   attribute ment_tsu83: string;
   attribute ment_tsu83 of DEF_ARCH : architecture is " F_FM0_WDATA[5]->CLK_BASE=0.494";
   attribute ment_tsu84: string;
   attribute ment_tsu84 of DEF_ARCH : architecture is " F_FM0_WDATA[6]->CLK_BASE=0.375";
   attribute ment_tsu85: string;
   attribute ment_tsu85 of DEF_ARCH : architecture is " F_FM0_WDATA[7]->CLK_BASE=0.367";
   attribute ment_tsu86: string;
   attribute ment_tsu86 of DEF_ARCH : architecture is " F_FM0_WDATA[8]->CLK_BASE=0.371";
   attribute ment_tsu87: string;
   attribute ment_tsu87 of DEF_ARCH : architecture is " F_FM0_WDATA[9]->CLK_BASE=0.360";
   attribute ment_tsu88: string;
   attribute ment_tsu88 of DEF_ARCH : architecture is " F_FM0_WRITE->CLK_BASE=0.562";
   attribute ment_tsu89: string;
   attribute ment_tsu89 of DEF_ARCH : architecture is " F_HM0_RDATA[0]->CLK_BASE=0.353";
   attribute ment_tsu90: string;
   attribute ment_tsu90 of DEF_ARCH : architecture is " F_HM0_RDATA[10]->CLK_BASE=0.365";
   attribute ment_tsu91: string;
   attribute ment_tsu91 of DEF_ARCH : architecture is " F_HM0_RDATA[11]->CLK_BASE=0.388";
   attribute ment_tsu92: string;
   attribute ment_tsu92 of DEF_ARCH : architecture is " F_HM0_RDATA[12]->CLK_BASE=0.516";
   attribute ment_tsu93: string;
   attribute ment_tsu93 of DEF_ARCH : architecture is " F_HM0_RDATA[13]->CLK_BASE=0.308";
   attribute ment_tsu94: string;
   attribute ment_tsu94 of DEF_ARCH : architecture is " F_HM0_RDATA[14]->CLK_BASE=0.339";
   attribute ment_tsu95: string;
   attribute ment_tsu95 of DEF_ARCH : architecture is " F_HM0_RDATA[15]->CLK_BASE=0.351";
   attribute ment_tsu96: string;
   attribute ment_tsu96 of DEF_ARCH : architecture is " F_HM0_RDATA[16]->CLK_BASE=0.405";
   attribute ment_tsu97: string;
   attribute ment_tsu97 of DEF_ARCH : architecture is " F_HM0_RDATA[17]->CLK_BASE=0.461";
   attribute ment_tsu98: string;
   attribute ment_tsu98 of DEF_ARCH : architecture is " F_HM0_RDATA[18]->CLK_BASE=0.460";
   attribute ment_tsu99: string;
   attribute ment_tsu99 of DEF_ARCH : architecture is " F_HM0_RDATA[19]->CLK_BASE=0.306";
   attribute ment_tsu100: string;
   attribute ment_tsu100 of DEF_ARCH : architecture is " F_HM0_RDATA[1]->CLK_BASE=0.440";
   attribute ment_tsu101: string;
   attribute ment_tsu101 of DEF_ARCH : architecture is " F_HM0_RDATA[20]->CLK_BASE=0.329";
   attribute ment_tsu102: string;
   attribute ment_tsu102 of DEF_ARCH : architecture is " F_HM0_RDATA[21]->CLK_BASE=0.400";
   attribute ment_tsu103: string;
   attribute ment_tsu103 of DEF_ARCH : architecture is " F_HM0_RDATA[22]->CLK_BASE=0.418";
   attribute ment_tsu104: string;
   attribute ment_tsu104 of DEF_ARCH : architecture is " F_HM0_RDATA[23]->CLK_BASE=0.427";
   attribute ment_tsu105: string;
   attribute ment_tsu105 of DEF_ARCH : architecture is " F_HM0_RDATA[24]->CLK_BASE=0.338";
   attribute ment_tsu106: string;
   attribute ment_tsu106 of DEF_ARCH : architecture is " F_HM0_RDATA[25]->CLK_BASE=0.381";
   attribute ment_tsu107: string;
   attribute ment_tsu107 of DEF_ARCH : architecture is " F_HM0_RDATA[26]->CLK_BASE=0.331";
   attribute ment_tsu108: string;
   attribute ment_tsu108 of DEF_ARCH : architecture is " F_HM0_RDATA[27]->CLK_BASE=0.369";
   attribute ment_tsu109: string;
   attribute ment_tsu109 of DEF_ARCH : architecture is " F_HM0_RDATA[28]->CLK_BASE=0.429";
   attribute ment_tsu110: string;
   attribute ment_tsu110 of DEF_ARCH : architecture is " F_HM0_RDATA[29]->CLK_BASE=0.425";
   attribute ment_tsu111: string;
   attribute ment_tsu111 of DEF_ARCH : architecture is " F_HM0_RDATA[2]->CLK_BASE=0.336";
   attribute ment_tsu112: string;
   attribute ment_tsu112 of DEF_ARCH : architecture is " F_HM0_RDATA[30]->CLK_BASE=0.414";
   attribute ment_tsu113: string;
   attribute ment_tsu113 of DEF_ARCH : architecture is " F_HM0_RDATA[31]->CLK_BASE=0.435";
   attribute ment_tsu114: string;
   attribute ment_tsu114 of DEF_ARCH : architecture is " F_HM0_RDATA[3]->CLK_BASE=0.346";
   attribute ment_tsu115: string;
   attribute ment_tsu115 of DEF_ARCH : architecture is " F_HM0_RDATA[4]->CLK_BASE=0.372";
   attribute ment_tsu116: string;
   attribute ment_tsu116 of DEF_ARCH : architecture is " F_HM0_RDATA[5]->CLK_BASE=0.428";
   attribute ment_tsu117: string;
   attribute ment_tsu117 of DEF_ARCH : architecture is " F_HM0_RDATA[6]->CLK_BASE=0.375";
   attribute ment_tsu118: string;
   attribute ment_tsu118 of DEF_ARCH : architecture is " F_HM0_RDATA[7]->CLK_BASE=0.353";
   attribute ment_tsu119: string;
   attribute ment_tsu119 of DEF_ARCH : architecture is " F_HM0_RDATA[8]->CLK_BASE=0.369";
   attribute ment_tsu120: string;
   attribute ment_tsu120 of DEF_ARCH : architecture is " F_HM0_RDATA[9]->CLK_BASE=0.348";
   attribute ment_tsu121: string;
   attribute ment_tsu121 of DEF_ARCH : architecture is " F_HM0_READY->CLK_BASE=1.479";
   attribute ment_tsu122: string;
   attribute ment_tsu122 of DEF_ARCH : architecture is " F_HM0_RESP->CLK_BASE=0.708";
   attribute ment_tsu123: string;
   attribute ment_tsu123 of DEF_ARCH : architecture is " I2C0_SDA_F2H_SCP->I2C0_SCL_F2H_SCP=0.195";
   attribute ment_tsu124: string;
   attribute ment_tsu124 of DEF_ARCH : architecture is " I2C1_SDA_F2H_SCP->I2C1_SCL_F2H_SCP=0.276";
   attribute ment_tsu125: string;
   attribute ment_tsu125 of DEF_ARCH : architecture is " MGPIO0A_F2H_GPIN->CLK_BASE=0.619";
   attribute ment_tsu126: string;
   attribute ment_tsu126 of DEF_ARCH : architecture is " MGPIO10A_F2H_GPIN->CLK_BASE=0.477";
   attribute ment_tsu127: string;
   attribute ment_tsu127 of DEF_ARCH : architecture is " MGPIO11A_F2H_GPIN->CLK_BASE=0.557";
   attribute ment_tsu128: string;
   attribute ment_tsu128 of DEF_ARCH : architecture is " MGPIO11B_F2H_GPIN->CLK_BASE=0.596";
   attribute ment_tsu129: string;
   attribute ment_tsu129 of DEF_ARCH : architecture is " MGPIO12A_F2H_GPIN->CLK_BASE=0.639";
   attribute ment_tsu130: string;
   attribute ment_tsu130 of DEF_ARCH : architecture is " MGPIO13A_F2H_GPIN->CLK_BASE=0.562";
   attribute ment_tsu131: string;
   attribute ment_tsu131 of DEF_ARCH : architecture is " MGPIO14A_F2H_GPIN->CLK_BASE=0.633";
   attribute ment_tsu132: string;
   attribute ment_tsu132 of DEF_ARCH : architecture is " MGPIO15A_F2H_GPIN->CLK_BASE=0.665";
   attribute ment_tsu133: string;
   attribute ment_tsu133 of DEF_ARCH : architecture is " MGPIO16A_F2H_GPIN->CLK_BASE=0.541";
   attribute ment_tsu134: string;
   attribute ment_tsu134 of DEF_ARCH : architecture is " MGPIO17B_F2H_GPIN->CLK_BASE=0.555";
   attribute ment_tsu135: string;
   attribute ment_tsu135 of DEF_ARCH : architecture is " MGPIO18B_F2H_GPIN->CLK_BASE=0.687";
   attribute ment_tsu136: string;
   attribute ment_tsu136 of DEF_ARCH : architecture is " MGPIO19B_F2H_GPIN->CLK_BASE=0.629";
   attribute ment_tsu137: string;
   attribute ment_tsu137 of DEF_ARCH : architecture is " MGPIO1A_F2H_GPIN->CLK_BASE=0.574";
   attribute ment_tsu138: string;
   attribute ment_tsu138 of DEF_ARCH : architecture is " MGPIO20B_F2H_GPIN->CLK_BASE=0.710";
   attribute ment_tsu139: string;
   attribute ment_tsu139 of DEF_ARCH : architecture is " MGPIO21B_F2H_GPIN->CLK_BASE=0.591";
   attribute ment_tsu140: string;
   attribute ment_tsu140 of DEF_ARCH : architecture is " MGPIO22B_F2H_GPIN->CLK_BASE=0.658";
   attribute ment_tsu141: string;
   attribute ment_tsu141 of DEF_ARCH : architecture is " MGPIO24B_F2H_GPIN->CLK_BASE=0.562";
   attribute ment_tsu142: string;
   attribute ment_tsu142 of DEF_ARCH : architecture is " MGPIO25B_F2H_GPIN->CLK_BASE=0.668";
   attribute ment_tsu143: string;
   attribute ment_tsu143 of DEF_ARCH : architecture is " MGPIO26B_F2H_GPIN->CLK_BASE=0.696";
   attribute ment_tsu144: string;
   attribute ment_tsu144 of DEF_ARCH : architecture is " MGPIO27B_F2H_GPIN->CLK_BASE=0.648";
   attribute ment_tsu145: string;
   attribute ment_tsu145 of DEF_ARCH : architecture is " MGPIO28B_F2H_GPIN->CLK_BASE=0.724";
   attribute ment_tsu146: string;
   attribute ment_tsu146 of DEF_ARCH : architecture is " MGPIO29B_F2H_GPIN->CLK_BASE=0.933";
   attribute ment_tsu147: string;
   attribute ment_tsu147 of DEF_ARCH : architecture is " MGPIO2A_F2H_GPIN->CLK_BASE=0.659";
   attribute ment_tsu148: string;
   attribute ment_tsu148 of DEF_ARCH : architecture is " MGPIO30B_F2H_GPIN->CLK_BASE=0.652";
   attribute ment_tsu149: string;
   attribute ment_tsu149 of DEF_ARCH : architecture is " MGPIO31B_F2H_GPIN->CLK_BASE=0.822";
   attribute ment_tsu150: string;
   attribute ment_tsu150 of DEF_ARCH : architecture is " MGPIO3A_F2H_GPIN->CLK_BASE=0.541";
   attribute ment_tsu151: string;
   attribute ment_tsu151 of DEF_ARCH : architecture is " MGPIO4A_F2H_GPIN->CLK_BASE=0.776";
   attribute ment_tsu152: string;
   attribute ment_tsu152 of DEF_ARCH : architecture is " MGPIO5A_F2H_GPIN->CLK_BASE=0.698";
   attribute ment_tsu153: string;
   attribute ment_tsu153 of DEF_ARCH : architecture is " MGPIO6A_F2H_GPIN->CLK_BASE=0.586";
   attribute ment_tsu154: string;
   attribute ment_tsu154 of DEF_ARCH : architecture is " MGPIO7A_F2H_GPIN->CLK_BASE=0.633";
   attribute ment_tsu155: string;
   attribute ment_tsu155 of DEF_ARCH : architecture is " MGPIO8A_F2H_GPIN->CLK_BASE=0.697";
   attribute ment_tsu156: string;
   attribute ment_tsu156 of DEF_ARCH : architecture is " MGPIO9A_F2H_GPIN->CLK_BASE=0.481";
   attribute ment_tsu157: string;
   attribute ment_tsu157 of DEF_ARCH : architecture is " MMUART0_CTS_F2H_SCP->CLK_BASE=1.134";
   attribute ment_tsu158: string;
   attribute ment_tsu158 of DEF_ARCH : architecture is " MMUART0_DCD_F2H_SCP->CLK_BASE=1.207";
   attribute ment_tsu159: string;
   attribute ment_tsu159 of DEF_ARCH : architecture is " MMUART0_DSR_F2H_SCP->CLK_BASE=1.158";
   attribute ment_tsu160: string;
   attribute ment_tsu160 of DEF_ARCH : architecture is " MMUART0_RI_F2H_SCP->CLK_BASE=0.821";
   attribute ment_tsu161: string;
   attribute ment_tsu161 of DEF_ARCH : architecture is " MMUART0_RXD_F2H_SCP->CLK_BASE=0.939";
   attribute ment_tsu162: string;
   attribute ment_tsu162 of DEF_ARCH : architecture is " MMUART0_SCK_F2H_SCP->CLK_BASE=1.070";
   attribute ment_tsu163: string;
   attribute ment_tsu163 of DEF_ARCH : architecture is " MMUART0_TXD_F2H_SCP->CLK_BASE=1.203";
   attribute ment_tsu164: string;
   attribute ment_tsu164 of DEF_ARCH : architecture is " MMUART1_CTS_F2H_SCP->CLK_BASE=1.051";
   attribute ment_tsu165: string;
   attribute ment_tsu165 of DEF_ARCH : architecture is " MMUART1_DCD_F2H_SCP->CLK_BASE=0.924";
   attribute ment_tsu166: string;
   attribute ment_tsu166 of DEF_ARCH : architecture is " MMUART1_DSR_F2H_SCP->CLK_BASE=1.010";
   attribute ment_tsu167: string;
   attribute ment_tsu167 of DEF_ARCH : architecture is " MMUART1_RI_F2H_SCP->CLK_BASE=0.814";
   attribute ment_tsu168: string;
   attribute ment_tsu168 of DEF_ARCH : architecture is " MMUART1_RXD_F2H_SCP->CLK_BASE=1.174";
   attribute ment_tsu169: string;
   attribute ment_tsu169 of DEF_ARCH : architecture is " MMUART1_SCK_F2H_SCP->CLK_BASE=0.802";
   attribute ment_tsu170: string;
   attribute ment_tsu170 of DEF_ARCH : architecture is " MMUART1_TXD_F2H_SCP->CLK_BASE=1.053";
   attribute ment_tsu171: string;
   attribute ment_tsu171 of DEF_ARCH : architecture is " SMBALERT_NI0->I2C0_SCL_F2H_SCP=-0.411";
   attribute ment_tsu172: string;
   attribute ment_tsu172 of DEF_ARCH : architecture is " SMBALERT_NI1->I2C1_SCL_F2H_SCP=-0.115";
   attribute ment_tsu173: string;
   attribute ment_tsu173 of DEF_ARCH : architecture is " SMBSUS_NI0->I2C0_SCL_F2H_SCP=-0.369";
   attribute ment_tsu174: string;
   attribute ment_tsu174 of DEF_ARCH : architecture is " SMBSUS_NI1->I2C1_SCL_F2H_SCP=-0.156";
   attribute ment_tsu175: string;
   attribute ment_tsu175 of DEF_ARCH : architecture is " SPI0_SDI_F2H_SCP->SPI0_CLK_IN=1.351";
   attribute ment_tsu176: string;
   attribute ment_tsu176 of DEF_ARCH : architecture is " SPI1_SDI_F2H_SCP->SPI1_CLK_IN=1.194";
   attribute ment_tco0: string;
   attribute ment_tco0 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_A=3.406";
   attribute ment_tco1: string;
   attribute ment_tco1 of DEF_ARCH : architecture is " CLK_BASE->CAN_RXBUS_MGPIO3A_H2F_B=3.430";
   attribute ment_tco2: string;
   attribute ment_tco2 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_A=3.332";
   attribute ment_tco3: string;
   attribute ment_tco3 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_MGPIO2A_H2F_B=3.416";
   attribute ment_tco4: string;
   attribute ment_tco4 of DEF_ARCH : architecture is " CLK_BASE->CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT=3.805";
   attribute ment_tco5: string;
   attribute ment_tco5 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_A=3.405";
   attribute ment_tco6: string;
   attribute ment_tco6 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_MGPIO4A_H2F_B=3.306";
   attribute ment_tco7: string;
   attribute ment_tco7 of DEF_ARCH : architecture is " CLK_BASE->CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT=3.712";
   attribute ment_tco8: string;
   attribute ment_tco8 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[0]=4.256";
   attribute ment_tco9: string;
   attribute ment_tco9 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[10]=4.211";
   attribute ment_tco10: string;
   attribute ment_tco10 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[11]=4.111";
   attribute ment_tco11: string;
   attribute ment_tco11 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[12]=4.281";
   attribute ment_tco12: string;
   attribute ment_tco12 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[13]=4.282";
   attribute ment_tco13: string;
   attribute ment_tco13 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[14]=4.165";
   attribute ment_tco14: string;
   attribute ment_tco14 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[15]=4.116";
   attribute ment_tco15: string;
   attribute ment_tco15 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[16]=4.196";
   attribute ment_tco16: string;
   attribute ment_tco16 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[17]=4.200";
   attribute ment_tco17: string;
   attribute ment_tco17 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[18]=4.173";
   attribute ment_tco18: string;
   attribute ment_tco18 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[19]=4.202";
   attribute ment_tco19: string;
   attribute ment_tco19 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[1]=4.144";
   attribute ment_tco20: string;
   attribute ment_tco20 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[20]=4.240";
   attribute ment_tco21: string;
   attribute ment_tco21 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[21]=4.233";
   attribute ment_tco22: string;
   attribute ment_tco22 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[22]=4.200";
   attribute ment_tco23: string;
   attribute ment_tco23 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[23]=4.190";
   attribute ment_tco24: string;
   attribute ment_tco24 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[24]=4.228";
   attribute ment_tco25: string;
   attribute ment_tco25 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[25]=4.219";
   attribute ment_tco26: string;
   attribute ment_tco26 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[26]=4.182";
   attribute ment_tco27: string;
   attribute ment_tco27 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[27]=4.271";
   attribute ment_tco28: string;
   attribute ment_tco28 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[28]=4.233";
   attribute ment_tco29: string;
   attribute ment_tco29 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[29]=4.248";
   attribute ment_tco30: string;
   attribute ment_tco30 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[2]=4.240";
   attribute ment_tco31: string;
   attribute ment_tco31 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[30]=4.150";
   attribute ment_tco32: string;
   attribute ment_tco32 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[31]=4.166";
   attribute ment_tco33: string;
   attribute ment_tco33 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[3]=4.263";
   attribute ment_tco34: string;
   attribute ment_tco34 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[4]=4.196";
   attribute ment_tco35: string;
   attribute ment_tco35 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[5]=4.117";
   attribute ment_tco36: string;
   attribute ment_tco36 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[6]=4.080";
   attribute ment_tco37: string;
   attribute ment_tco37 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[7]=4.125";
   attribute ment_tco38: string;
   attribute ment_tco38 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[8]=4.202";
   attribute ment_tco39: string;
   attribute ment_tco39 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RDATA[9]=4.098";
   attribute ment_tco40: string;
   attribute ment_tco40 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_READYOUT=3.920";
   attribute ment_tco41: string;
   attribute ment_tco41 of DEF_ARCH : architecture is " CLK_BASE->F_FM0_RESP=3.932";
   attribute ment_tco42: string;
   attribute ment_tco42 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[0]=3.432";
   attribute ment_tco43: string;
   attribute ment_tco43 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[10]=3.216";
   attribute ment_tco44: string;
   attribute ment_tco44 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[11]=3.231";
   attribute ment_tco45: string;
   attribute ment_tco45 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[12]=3.172";
   attribute ment_tco46: string;
   attribute ment_tco46 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[13]=3.213";
   attribute ment_tco47: string;
   attribute ment_tco47 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[14]=3.180";
   attribute ment_tco48: string;
   attribute ment_tco48 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[15]=3.206";
   attribute ment_tco49: string;
   attribute ment_tco49 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[16]=3.223";
   attribute ment_tco50: string;
   attribute ment_tco50 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[17]=3.219";
   attribute ment_tco51: string;
   attribute ment_tco51 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[18]=3.207";
   attribute ment_tco52: string;
   attribute ment_tco52 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[19]=3.195";
   attribute ment_tco53: string;
   attribute ment_tco53 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[1]=3.474";
   attribute ment_tco54: string;
   attribute ment_tco54 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[20]=3.188";
   attribute ment_tco55: string;
   attribute ment_tco55 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[21]=3.191";
   attribute ment_tco56: string;
   attribute ment_tco56 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[22]=3.213";
   attribute ment_tco57: string;
   attribute ment_tco57 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[23]=3.246";
   attribute ment_tco58: string;
   attribute ment_tco58 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[24]=3.163";
   attribute ment_tco59: string;
   attribute ment_tco59 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[25]=3.197";
   attribute ment_tco60: string;
   attribute ment_tco60 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[26]=3.239";
   attribute ment_tco61: string;
   attribute ment_tco61 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[27]=3.195";
   attribute ment_tco62: string;
   attribute ment_tco62 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[28]=3.230";
   attribute ment_tco63: string;
   attribute ment_tco63 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[29]=3.161";
   attribute ment_tco64: string;
   attribute ment_tco64 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[2]=3.235";
   attribute ment_tco65: string;
   attribute ment_tco65 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[30]=3.194";
   attribute ment_tco66: string;
   attribute ment_tco66 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[31]=3.230";
   attribute ment_tco67: string;
   attribute ment_tco67 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[3]=3.200";
   attribute ment_tco68: string;
   attribute ment_tco68 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[4]=3.205";
   attribute ment_tco69: string;
   attribute ment_tco69 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[5]=3.222";
   attribute ment_tco70: string;
   attribute ment_tco70 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[6]=3.203";
   attribute ment_tco71: string;
   attribute ment_tco71 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[7]=3.191";
   attribute ment_tco72: string;
   attribute ment_tco72 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[8]=3.244";
   attribute ment_tco73: string;
   attribute ment_tco73 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_ADDR[9]=3.191";
   attribute ment_tco74: string;
   attribute ment_tco74 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SEL=3.323";
   attribute ment_tco75: string;
   attribute ment_tco75 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SIZE[0]=3.310";
   attribute ment_tco76: string;
   attribute ment_tco76 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_SIZE[1]=3.357";
   attribute ment_tco77: string;
   attribute ment_tco77 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_TRANS1=3.228";
   attribute ment_tco78: string;
   attribute ment_tco78 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[0]=3.170";
   attribute ment_tco79: string;
   attribute ment_tco79 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[10]=3.311";
   attribute ment_tco80: string;
   attribute ment_tco80 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[11]=3.361";
   attribute ment_tco81: string;
   attribute ment_tco81 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[12]=3.298";
   attribute ment_tco82: string;
   attribute ment_tco82 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[13]=3.446";
   attribute ment_tco83: string;
   attribute ment_tco83 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[14]=3.230";
   attribute ment_tco84: string;
   attribute ment_tco84 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[15]=3.356";
   attribute ment_tco85: string;
   attribute ment_tco85 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[16]=3.330";
   attribute ment_tco86: string;
   attribute ment_tco86 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[17]=3.371";
   attribute ment_tco87: string;
   attribute ment_tco87 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[18]=3.302";
   attribute ment_tco88: string;
   attribute ment_tco88 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[19]=3.431";
   attribute ment_tco89: string;
   attribute ment_tco89 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[1]=3.176";
   attribute ment_tco90: string;
   attribute ment_tco90 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[20]=3.304";
   attribute ment_tco91: string;
   attribute ment_tco91 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[21]=3.422";
   attribute ment_tco92: string;
   attribute ment_tco92 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[22]=3.386";
   attribute ment_tco93: string;
   attribute ment_tco93 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[23]=3.099";
   attribute ment_tco94: string;
   attribute ment_tco94 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[24]=3.293";
   attribute ment_tco95: string;
   attribute ment_tco95 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[25]=3.447";
   attribute ment_tco96: string;
   attribute ment_tco96 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[26]=3.480";
   attribute ment_tco97: string;
   attribute ment_tco97 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[27]=3.444";
   attribute ment_tco98: string;
   attribute ment_tco98 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[28]=3.418";
   attribute ment_tco99: string;
   attribute ment_tco99 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[29]=3.478";
   attribute ment_tco100: string;
   attribute ment_tco100 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[2]=3.256";
   attribute ment_tco101: string;
   attribute ment_tco101 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[30]=3.531";
   attribute ment_tco102: string;
   attribute ment_tco102 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[31]=3.483";
   attribute ment_tco103: string;
   attribute ment_tco103 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[3]=3.114";
   attribute ment_tco104: string;
   attribute ment_tco104 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[4]=3.310";
   attribute ment_tco105: string;
   attribute ment_tco105 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[5]=3.299";
   attribute ment_tco106: string;
   attribute ment_tco106 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[6]=3.386";
   attribute ment_tco107: string;
   attribute ment_tco107 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[7]=3.393";
   attribute ment_tco108: string;
   attribute ment_tco108 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[8]=3.399";
   attribute ment_tco109: string;
   attribute ment_tco109 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WDATA[9]=3.388";
   attribute ment_tco110: string;
   attribute ment_tco110 of DEF_ARCH : architecture is " CLK_BASE->F_HM0_WRITE=3.628";
   attribute ment_tco111: string;
   attribute ment_tco111 of DEF_ARCH : architecture is " CLK_BASE->H2FCALIB=3.101";
   attribute ment_tco112: string;
   attribute ment_tco112 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_MGPIO31B_H2F_B=3.461";
   attribute ment_tco113: string;
   attribute ment_tco113 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SCL_USBC_DATA1_MGPIO31B_OE=3.462";
   attribute ment_tco114: string;
   attribute ment_tco114 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_A=3.507";
   attribute ment_tco115: string;
   attribute ment_tco115 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_MGPIO30B_H2F_B=3.405";
   attribute ment_tco116: string;
   attribute ment_tco116 of DEF_ARCH : architecture is " CLK_BASE->I2C0_SDA_USBC_DATA0_MGPIO30B_OE=2.892";
   attribute ment_tco117: string;
   attribute ment_tco117 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_MGPIO1A_H2F_B=3.412";
   attribute ment_tco118: string;
   attribute ment_tco118 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SCL_USBA_DATA4_MGPIO1A_OE=3.434";
   attribute ment_tco119: string;
   attribute ment_tco119 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_A=3.354";
   attribute ment_tco120: string;
   attribute ment_tco120 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_MGPIO0A_H2F_B=3.505";
   attribute ment_tco121: string;
   attribute ment_tco121 of DEF_ARCH : architecture is " CLK_BASE->I2C1_SDA_USBA_DATA3_MGPIO0A_OE=3.338";
   attribute ment_tco122: string;
   attribute ment_tco122 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OE=2.796";
   attribute ment_tco123: string;
   attribute ment_tco123 of DEF_ARCH : architecture is " CLK_BASE->MGPIO25A_OUT=2.714";
   attribute ment_tco124: string;
   attribute ment_tco124 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OE=2.752";
   attribute ment_tco125: string;
   attribute ment_tco125 of DEF_ARCH : architecture is " CLK_BASE->MGPIO26A_OUT=2.837";
   attribute ment_tco126: string;
   attribute ment_tco126 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_A=3.371";
   attribute ment_tco127: string;
   attribute ment_tco127 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_CTS_MGPIO19B_H2F_B=3.512";
   attribute ment_tco128: string;
   attribute ment_tco128 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_A=3.236";
   attribute ment_tco129: string;
   attribute ment_tco129 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DCD_MGPIO22B_H2F_B=3.402";
   attribute ment_tco130: string;
   attribute ment_tco130 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_A=3.263";
   attribute ment_tco131: string;
   attribute ment_tco131 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DSR_MGPIO20B_H2F_B=3.450";
   attribute ment_tco132: string;
   attribute ment_tco132 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_A=3.241";
   attribute ment_tco133: string;
   attribute ment_tco133 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_MGPIO18B_H2F_B=3.368";
   attribute ment_tco134: string;
   attribute ment_tco134 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT=2.834";
   attribute ment_tco135: string;
   attribute ment_tco135 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_A=3.459";
   attribute ment_tco136: string;
   attribute ment_tco136 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RI_MGPIO21B_H2F_B=3.419";
   attribute ment_tco137: string;
   attribute ment_tco137 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_A=3.450";
   attribute ment_tco138: string;
   attribute ment_tco138 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_MGPIO17B_H2F_B=3.406";
   attribute ment_tco139: string;
   attribute ment_tco139 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT=2.950";
   attribute ment_tco140: string;
   attribute ment_tco140 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_A=3.514";
   attribute ment_tco141: string;
   attribute ment_tco141 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_RXD_MGPIO28B_H2F_B=3.434";
   attribute ment_tco142: string;
   attribute ment_tco142 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_A=3.289";
   attribute ment_tco143: string;
   attribute ment_tco143 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_MGPIO29B_H2F_B=3.407";
   attribute ment_tco144: string;
   attribute ment_tco144 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OE=3.181";
   attribute ment_tco145: string;
   attribute ment_tco145 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_SCK_USBC_NXT_MGPIO29B_OUT=2.738";
   attribute ment_tco146: string;
   attribute ment_tco146 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_A=3.507";
   attribute ment_tco147: string;
   attribute ment_tco147 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_MGPIO27B_H2F_B=3.404";
   attribute ment_tco148: string;
   attribute ment_tco148 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OE=3.439";
   attribute ment_tco149: string;
   attribute ment_tco149 of DEF_ARCH : architecture is " CLK_BASE->MMUART0_TXD_USBC_DIR_MGPIO27B_OUT=2.938";
   attribute ment_tco150: string;
   attribute ment_tco150 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_H2F_A=3.359";
   attribute ment_tco151: string;
   attribute ment_tco151 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_DTR_MGPIO12B_OUT=3.084";
   attribute ment_tco152: string;
   attribute ment_tco152 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_A=3.350";
   attribute ment_tco153: string;
   attribute ment_tco153 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_H2F_B=3.401";
   attribute ment_tco154: string;
   attribute ment_tco154 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RTS_MGPIO11B_OUT=3.048";
   attribute ment_tco155: string;
   attribute ment_tco155 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_A=3.474";
   attribute ment_tco156: string;
   attribute ment_tco156 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_RXD_MGPIO26B_H2F_B=3.183";
   attribute ment_tco157: string;
   attribute ment_tco157 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_A=3.283";
   attribute ment_tco158: string;
   attribute ment_tco158 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_MGPIO25B_H2F_B=3.474";
   attribute ment_tco159: string;
   attribute ment_tco159 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OE=3.652";
   attribute ment_tco160: string;
   attribute ment_tco160 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT=2.702";
   attribute ment_tco161: string;
   attribute ment_tco161 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_A=3.431";
   attribute ment_tco162: string;
   attribute ment_tco162 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_MGPIO24B_H2F_B=4.408";
   attribute ment_tco163: string;
   attribute ment_tco163 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OE=3.431";
   attribute ment_tco164: string;
   attribute ment_tco164 of DEF_ARCH : architecture is " CLK_BASE->MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT=3.287";
   attribute ment_tco165: string;
   attribute ment_tco165 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE=3.917";
   attribute ment_tco166: string;
   attribute ment_tco166 of DEF_ARCH : architecture is " CLK_BASE->RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT=4.161";
   attribute ment_tco167: string;
   attribute ment_tco167 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_A=3.513";
   attribute ment_tco168: string;
   attribute ment_tco168 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDI_MGPIO5A_H2F_B=3.511";
   attribute ment_tco169: string;
   attribute ment_tco169 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_A=3.581";
   attribute ment_tco170: string;
   attribute ment_tco170 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_MGPIO6A_H2F_B=3.494";
   attribute ment_tco171: string;
   attribute ment_tco171 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OE=5.005";
   attribute ment_tco172: string;
   attribute ment_tco172 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SDO_USBA_STP_MGPIO6A_OUT=5.220";
   attribute ment_tco173: string;
   attribute ment_tco173 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_A=3.367";
   attribute ment_tco174: string;
   attribute ment_tco174 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS0_MGPIO7A_H2F_B=3.467";
   attribute ment_tco175: string;
   attribute ment_tco175 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_A=3.499";
   attribute ment_tco176: string;
   attribute ment_tco176 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS1_MGPIO8A_H2F_B=3.524";
   attribute ment_tco177: string;
   attribute ment_tco177 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_A=3.334";
   attribute ment_tco178: string;
   attribute ment_tco178 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS2_MGPIO9A_H2F_B=3.361";
   attribute ment_tco179: string;
   attribute ment_tco179 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_A=3.390";
   attribute ment_tco180: string;
   attribute ment_tco180 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS3_MGPIO10A_H2F_B=3.446";
   attribute ment_tco181: string;
   attribute ment_tco181 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS4_MGPIO19A_H2F_A=3.529";
   attribute ment_tco182: string;
   attribute ment_tco182 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS5_MGPIO20A_H2F_A=3.217";
   attribute ment_tco183: string;
   attribute ment_tco183 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS6_MGPIO21A_H2F_A=3.402";
   attribute ment_tco184: string;
   attribute ment_tco184 of DEF_ARCH : architecture is " CLK_BASE->SPI0_SS7_MGPIO22A_H2F_A=3.630";
   attribute ment_tco185: string;
   attribute ment_tco185 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_A=3.584";
   attribute ment_tco186: string;
   attribute ment_tco186 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDI_MGPIO11A_H2F_B=3.903";
   attribute ment_tco187: string;
   attribute ment_tco187 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_A=3.223";
   attribute ment_tco188: string;
   attribute ment_tco188 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_H2F_B=3.372";
   attribute ment_tco189: string;
   attribute ment_tco189 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OE=5.380";
   attribute ment_tco190: string;
   attribute ment_tco190 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SDO_MGPIO12A_OUT=5.553";
   attribute ment_tco191: string;
   attribute ment_tco191 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_A=3.832";
   attribute ment_tco192: string;
   attribute ment_tco192 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS0_MGPIO13A_H2F_B=4.024";
   attribute ment_tco193: string;
   attribute ment_tco193 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_A=3.365";
   attribute ment_tco194: string;
   attribute ment_tco194 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS1_MGPIO14A_H2F_B=3.235";
   attribute ment_tco195: string;
   attribute ment_tco195 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_A=3.407";
   attribute ment_tco196: string;
   attribute ment_tco196 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS2_MGPIO15A_H2F_B=3.255";
   attribute ment_tco197: string;
   attribute ment_tco197 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_A=3.287";
   attribute ment_tco198: string;
   attribute ment_tco198 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS3_MGPIO16A_H2F_B=3.347";
   attribute ment_tco199: string;
   attribute ment_tco199 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS4_MGPIO17A_H2F_A=3.654";
   attribute ment_tco200: string;
   attribute ment_tco200 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS5_MGPIO18A_H2F_A=3.351";
   attribute ment_tco201: string;
   attribute ment_tco201 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS6_MGPIO23A_H2F_A=3.465";
   attribute ment_tco202: string;
   attribute ment_tco202 of DEF_ARCH : architecture is " CLK_BASE->SPI1_SS7_MGPIO24A_H2F_A=3.411";
   attribute black_box_pad : string;
   attribute black_box_pad of DEF_ARCH : architecture is "";

begin

end DEF_ARCH;
